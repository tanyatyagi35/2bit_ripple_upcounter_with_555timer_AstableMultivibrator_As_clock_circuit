* /home/tanyatyagi35/eSim-Workspace/ripplecounter_555timer_tanya/ripplecounter_555timer_tanya.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sat 08 Oct 2022 10:52:28 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U5  Net-_U3-Pad4_ Net-_U2-Pad6_ Net-_U4-Pad1_ Net-_U4-Pad2_ tanya_ripple_upcounter2		
U4  Net-_U4-Pad1_ Net-_U4-Pad2_ output1 output0 dac_bridge_2		
X1  Net-_X1-Pad1_ Net-_X1-Pad2_ Net-_C2-Pad2_ Net-_C1-Pad1_ Net-_U2-Pad2_ GND avsd_opamp		
X2  Net-_X1-Pad1_ Net-_X1-Pad2_ Net-_R2-Pad2_ Net-_C2-Pad2_ Net-_U2-Pad1_ GND avsd_opamp		
R1  Net-_R1-Pad1_ Net-_C1-Pad1_ 5k		
R2  Net-_C1-Pad1_ Net-_R2-Pad2_ 5k		
R3  Net-_R2-Pad2_ GND 5k		
R5  Net-_R1-Pad1_ Net-_Q1-Pad1_ 1k		
R4  Net-_Q1-Pad1_ Net-_C2-Pad2_ 2k		
C2  GND Net-_C2-Pad2_ 10u		
Q1  Net-_Q1-Pad1_ Net-_Q1-Pad2_ GND eSim_NPN		
C1  Net-_C1-Pad1_ GND 0.01u		
v1  Net-_R1-Pad1_ GND 5		
v5  Net-_X1-Pad1_ GND 1		
v4  GND Net-_X1-Pad2_ 1		
v6  Net-_U2-Pad3_ GND pulse		
U6  output1 plot_v1		
U7  output0 plot_v1		
U3  Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ Net-_U3-Pad4_ Net-_U1-Pad1_ tanya_srff		
U2  Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ adc_bridge_3		
U1  Net-_U1-Pad1_ Net-_Q1-Pad2_ dac_bridge_1		
scmode1  SKY130mode		

.end
